`timescale 1ns/1ps


`define SMEM_MAX 1024
`define RMEM_MAX 256
`define TRANSACTION_COUNT 100
`define DRIV_IF topif.ME_DRIVER.ME_driver_cb
`define MON_IF topif.ME_MONITOR.ME_monitor_cb
